--no modifications were made to the downcounter.vhd module for our lab4 design

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_downcounter is
end entity;


--apparently we dont need this for the demo 