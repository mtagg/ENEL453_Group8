library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4089	)	,
(	4078	)	,
(	4068	)	,
(	4057	)	,
(	4046	)	,
(	4036	)	,
(	4025	)	,
(	4015	)	,
(	4004	)	,
(	3994	)	,
(	3984	)	,
(	3973	)	,
(	3963	)	,
(	3953	)	,
(	3942	)	,
(	3932	)	,
(	3922	)	,
(	3912	)	,
(	3902	)	,
(	3891	)	,
(	3881	)	,
(	3871	)	,
(	3861	)	,
(	3851	)	,
(	3841	)	,
(	3831	)	,
(	3821	)	,
(	3811	)	,
(	3801	)	,
(	3791	)	,
(	3781	)	,
(	3772	)	,
(	3762	)	,
(	3752	)	,
(	3742	)	,
(	3732	)	,
(	3723	)	,
(	3713	)	,
(	3703	)	,
(	3694	)	,
(	3684	)	,
(	3674	)	,
(	3665	)	,
(	3655	)	,
(	3646	)	,
(	3636	)	,
(	3627	)	,
(	3617	)	,
(	3608	)	,
(	3599	)	,
(	3589	)	,
(	3580	)	,
(	3571	)	,
(	3561	)	,
(	3552	)	,
(	3543	)	,
(	3533	)	,
(	3524	)	,
(	3515	)	,
(	3506	)	,
(	3497	)	,
(	3488	)	,
(	3479	)	,
(	3470	)	,
(	3461	)	,
(	3452	)	,
(	3443	)	,
(	3434	)	,
(	3425	)	,
(	3416	)	,
(	3407	)	,
(	3398	)	,
(	3389	)	,
(	3380	)	,
(	3372	)	,
(	3363	)	,
(	3354	)	,
(	3345	)	,
(	3337	)	,
(	3328	)	,
(	3319	)	,
(	3311	)	,
(	3302	)	,
(	3293	)	,
(	3285	)	,
(	3276	)	,
(	3268	)	,
(	3259	)	,
(	3251	)	,
(	3242	)	,
(	3234	)	,
(	3226	)	,
(	3217	)	,
(	3209	)	,
(	3201	)	,
(	3192	)	,
(	3184	)	,
(	3176	)	,
(	3167	)	,
(	3159	)	,
(	3151	)	,
(	3143	)	,
(	3135	)	,
(	3127	)	,
(	3118	)	,
(	3110	)	,
(	3102	)	,
(	3094	)	,
(	3086	)	,
(	3078	)	,
(	3070	)	,
(	3062	)	,
(	3054	)	,
(	3046	)	,
(	3039	)	,
(	3031	)	,
(	3023	)	,
(	3015	)	,
(	3007	)	,
(	2999	)	,
(	2992	)	,
(	2984	)	,
(	2976	)	,
(	2969	)	,
(	2961	)	,
(	2953	)	,
(	2946	)	,
(	2938	)	,
(	2930	)	,
(	2923	)	,
(	2915	)	,
(	2908	)	,
(	2900	)	,
(	2893	)	,
(	2885	)	,
(	2878	)	,
(	2870	)	,
(	2863	)	,
(	2856	)	,
(	2848	)	,
(	2841	)	,
(	2834	)	,
(	2826	)	,
(	2819	)	,
(	2812	)	,
(	2805	)	,
(	2797	)	,
(	2790	)	,
(	2783	)	,
(	2776	)	,
(	2769	)	,
(	2762	)	,
(	2755	)	,
(	2748	)	,
(	2741	)	,
(	2734	)	,
(	2727	)	,
(	2720	)	,
(	2713	)	,
(	2706	)	,
(	2699	)	,
(	2692	)	,
(	2685	)	,
(	2678	)	,
(	2671	)	,
(	2664	)	,
(	2658	)	,
(	2651	)	,
(	2644	)	,
(	2637	)	,
(	2631	)	,
(	2624	)	,
(	2617	)	,
(	2611	)	,
(	2604	)	,
(	2597	)	,
(	2591	)	,
(	2584	)	,
(	2577	)	,
(	2571	)	,
(	2564	)	,
(	2558	)	,
(	2551	)	,
(	2545	)	,
(	2538	)	,
(	2532	)	,
(	2526	)	,
(	2519	)	,
(	2513	)	,
(	2506	)	,
(	2500	)	,
(	2494	)	,
(	2488	)	,
(	2481	)	,
(	2475	)	,
(	2469	)	,
(	2463	)	,
(	2456	)	,
(	2450	)	,
(	2444	)	,
(	2438	)	,
(	2432	)	,
(	2426	)	,
(	2419	)	,
(	2413	)	,
(	2407	)	,
(	2401	)	,
(	2395	)	,
(	2389	)	,
(	2383	)	,
(	2377	)	,
(	2371	)	,
(	2365	)	,
(	2359	)	,
(	2354	)	,
(	2348	)	,
(	2342	)	,
(	2336	)	,
(	2330	)	,
(	2324	)	,
(	2319	)	,
(	2313	)	,
(	2307	)	,
(	2301	)	,
(	2296	)	,
(	2290	)	,
(	2284	)	,
(	2279	)	,
(	2273	)	,
(	2267	)	,
(	2262	)	,
(	2256	)	,
(	2250	)	,
(	2245	)	,
(	2239	)	,
(	2234	)	,
(	2228	)	,
(	2223	)	,
(	2217	)	,
(	2212	)	,
(	2206	)	,
(	2201	)	,
(	2196	)	,
(	2190	)	,
(	2185	)	,
(	2180	)	,
(	2174	)	,
(	2169	)	,
(	2164	)	,
(	2158	)	,
(	2153	)	,
(	2148	)	,
(	2143	)	,
(	2137	)	,
(	2132	)	,
(	2127	)	,
(	2122	)	,
(	2117	)	,
(	2111	)	,
(	2106	)	,
(	2101	)	,
(	2096	)	,
(	2091	)	,
(	2086	)	,
(	2081	)	,
(	2076	)	,
(	2071	)	,
(	2066	)	,
(	2061	)	,
(	2056	)	,
(	2051	)	,
(	2046	)	,
(	2041	)	,
(	2036	)	,
(	2031	)	,
(	2027	)	,
(	2022	)	,
(	2017	)	,
(	2012	)	,
(	2007	)	,
(	2002	)	,
(	1998	)	,
(	1993	)	,
(	1988	)	,
(	1983	)	,
(	1979	)	,
(	1974	)	,
(	1969	)	,
(	1965	)	,
(	1960	)	,
(	1955	)	,
(	1951	)	,
(	1946	)	,
(	1942	)	,
(	1937	)	,
(	1932	)	,
(	1928	)	,
(	1923	)	,
(	1919	)	,
(	1914	)	,
(	1910	)	,
(	1905	)	,
(	1901	)	,
(	1897	)	,
(	1892	)	,
(	1888	)	,
(	1883	)	,
(	1879	)	,
(	1875	)	,
(	1870	)	,
(	1866	)	,
(	1862	)	,
(	1857	)	,
(	1853	)	,
(	1849	)	,
(	1844	)	,
(	1840	)	,
(	1836	)	,
(	1832	)	,
(	1828	)	,
(	1823	)	,
(	1819	)	,
(	1815	)	,
(	1811	)	,
(	1807	)	,
(	1803	)	,
(	1799	)	,
(	1794	)	,
(	1790	)	,
(	1786	)	,
(	1782	)	,
(	1778	)	,
(	1774	)	,
(	1770	)	,
(	1766	)	,
(	1762	)	,
(	1758	)	,
(	1754	)	,
(	1750	)	,
(	1746	)	,
(	1743	)	,
(	1739	)	,
(	1735	)	,
(	1731	)	,
(	1727	)	,
(	1723	)	,
(	1719	)	,
(	1716	)	,
(	1712	)	,
(	1708	)	,
(	1704	)	,
(	1700	)	,
(	1697	)	,
(	1693	)	,
(	1689	)	,
(	1686	)	,
(	1682	)	,
(	1678	)	,
(	1674	)	,
(	1671	)	,
(	1667	)	,
(	1664	)	,
(	1660	)	,
(	1656	)	,
(	1653	)	,
(	1649	)	,
(	1646	)	,
(	1642	)	,
(	1638	)	,
(	1635	)	,
(	1631	)	,
(	1628	)	,
(	1624	)	,
(	1621	)	,
(	1618	)	,
(	1614	)	,
(	1611	)	,
(	1607	)	,
(	1604	)	,
(	1600	)	,
(	1597	)	,
(	1594	)	,
(	1590	)	,
(	1587	)	,
(	1584	)	,
(	1580	)	,
(	1577	)	,
(	1574	)	,
(	1570	)	,
(	1567	)	,
(	1564	)	,
(	1560	)	,
(	1557	)	,
(	1554	)	,
(	1551	)	,
(	1548	)	,
(	1544	)	,
(	1541	)	,
(	1538	)	,
(	1535	)	,
(	1532	)	,
(	1529	)	,
(	1525	)	,
(	1522	)	,
(	1519	)	,
(	1516	)	,
(	1513	)	,
(	1510	)	,
(	1507	)	,
(	1504	)	,
(	1501	)	,
(	1498	)	,
(	1495	)	,
(	1492	)	,
(	1489	)	,
(	1486	)	,
(	1483	)	,
(	1480	)	,
(	1477	)	,
(	1474	)	,
(	1471	)	,
(	1468	)	,
(	1465	)	,
(	1462	)	,
(	1460	)	,
(	1457	)	,
(	1454	)	,
(	1451	)	,
(	1448	)	,
(	1445	)	,
(	1443	)	,
(	1440	)	,
(	1437	)	,
(	1434	)	,
(	1431	)	,
(	1429	)	,
(	1426	)	,
(	1423	)	,
(	1420	)	,
(	1418	)	,
(	1415	)	,
(	1412	)	,
(	1410	)	,
(	1407	)	,
(	1404	)	,
(	1402	)	,
(	1399	)	,
(	1396	)	,
(	1394	)	,
(	1391	)	,
(	1388	)	,
(	1386	)	,
(	1383	)	,
(	1381	)	,
(	1378	)	,
(	1376	)	,
(	1373	)	,
(	1371	)	,
(	1368	)	,
(	1366	)	,
(	1363	)	,
(	1361	)	,
(	1358	)	,
(	1356	)	,
(	1353	)	,
(	1351	)	,
(	1348	)	,
(	1346	)	,
(	1343	)	,
(	1341	)	,
(	1339	)	,
(	1336	)	,
(	1334	)	,
(	1331	)	,
(	1329	)	,
(	1327	)	,
(	1324	)	,
(	1322	)	,
(	1320	)	,
(	1317	)	,
(	1315	)	,
(	1313	)	,
(	1311	)	,
(	1308	)	,
(	1306	)	,
(	1304	)	,
(	1301	)	,
(	1299	)	,
(	1297	)	,
(	1295	)	,
(	1293	)	,
(	1290	)	,
(	1288	)	,
(	1286	)	,
(	1284	)	,
(	1282	)	,
(	1279	)	,
(	1277	)	,
(	1275	)	,
(	1273	)	,
(	1271	)	,
(	1269	)	,
(	1267	)	,
(	1265	)	,
(	1262	)	,
(	1260	)	,
(	1258	)	,
(	1256	)	,
(	1254	)	,
(	1252	)	,
(	1250	)	,
(	1248	)	,
(	1246	)	,
(	1244	)	,
(	1242	)	,
(	1240	)	,
(	1238	)	,
(	1236	)	,
(	1234	)	,
(	1232	)	,
(	1230	)	,
(	1228	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1221	)	,
(	1219	)	,
(	1217	)	,
(	1215	)	,
(	1213	)	,
(	1211	)	,
(	1209	)	,
(	1207	)	,
(	1206	)	,
(	1204	)	,
(	1202	)	,
(	1200	)	,
(	1198	)	,
(	1196	)	,
(	1195	)	,
(	1193	)	,
(	1191	)	,
(	1189	)	,
(	1188	)	,
(	1186	)	,
(	1184	)	,
(	1182	)	,
(	1181	)	,
(	1179	)	,
(	1177	)	,
(	1175	)	,
(	1174	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1167	)	,
(	1165	)	,
(	1164	)	,
(	1162	)	,
(	1160	)	,
(	1159	)	,
(	1157	)	,
(	1155	)	,
(	1154	)	,
(	1152	)	,
(	1151	)	,
(	1149	)	,
(	1147	)	,
(	1146	)	,
(	1144	)	,
(	1143	)	,
(	1141	)	,
(	1140	)	,
(	1138	)	,
(	1136	)	,
(	1135	)	,
(	1133	)	,
(	1132	)	,
(	1130	)	,
(	1129	)	,
(	1127	)	,
(	1126	)	,
(	1124	)	,
(	1123	)	,
(	1121	)	,
(	1120	)	,
(	1119	)	,
(	1117	)	,
(	1116	)	,
(	1114	)	,
(	1113	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1107	)	,
(	1106	)	,
(	1104	)	,
(	1103	)	,
(	1102	)	,
(	1100	)	,
(	1099	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1089	)	,
(	1088	)	,
(	1087	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1025	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	989	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	985	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	977	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	971	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	968	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	963	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	958	)	,
(	957	)	,
(	956	)	,
(	956	)	,
(	955	)	,
(	954	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	947	)	,
(	946	)	,
(	945	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	940	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	883	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	629	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	620	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	607	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	577	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	571	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	566	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	556	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	550	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	540	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	534	)	,
(	533	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	524	)	,
(	523	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	519	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	508	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	502	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	498	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	492	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	484	)	,
(	483	)	,
(	482	)	,
(	481	)	,
(	480	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	475	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	471	)	,
(	470	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	466	)	,
(	465	)	,
(	464	)	,
(	463	)	,
(	462	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	455	)	,
(	454	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	450	)	,
(	449	)	,
(	448	)	,
(	447	)	,
(	446	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	442	)	,
(	441	)	,
(	440	)	,
(	439	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	435	)	,
(	434	)	,
(	433	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	429	)	,
(	428	)	,
(	427	)	,
(	426	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	422	)	,
(	421	)	,
(	420	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	416	)	,
(	415	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	411	)	,
(	410	)	,
(	409	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	405	)	,
(	404	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	400	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	




);


end package LUT_pkg;
