library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

 package LUT_pkg is

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	3794	)	, -- array index 0 (voltage = "000000000000" or 0 mV), distance output 3794 (37.94 cm)
(	3792	)	, -- array index 1 (voltage = "000000000001" or 1 mV), distance output 3792 (37.92 cm)
(	3791	)	,
(	3790	)	,
(	3789	)	,
(	3787	)	, -- array index 5 (voltage = "000000000101" or 5 mV), distance output 3787 (37.87 cm)
(	3786	)	,
(	3785	)	,
(	3784	)	,
(	3783	)	,
(	3781	)	,
(	3780	)	,
(	3779	)	,
(	3778	)	,
(	3776	)	,
(	3775	)	,
(	3774	)	,
(	3773	)	,
(	3771	)	,
(	3770	)	,
(	3769	)	,
(	3768	)	,
(	3766	)	,
(	3765	)	,
(	3764	)	,
(	3763	)	,
(	3762	)	,
(	3760	)	,
(	3759	)	,
(	3758	)	,
(	3757	)	,
(	3755	)	,
(	3754	)	,
(	3753	)	,
(	3752	)	,
(	3750	)	,
(	3749	)	,
(	3748	)	,
(	3747	)	,
(	3745	)	,
(	3744	)	,
(	3743	)	,
(	3742	)	,
(	3741	)	,
(	3739	)	,
(	3738	)	,
(	3737	)	,
(	3736	)	,
(	3734	)	,
(	3733	)	,
(	3732	)	,
(	3731	)	,
(	3729	)	,
(	3728	)	,
(	3727	)	,
(	3726	)	,
(	3725	)	,
(	3723	)	,
(	3722	)	,
(	3721	)	,
(	3720	)	,
(	3718	)	,
(	3717	)	,
(	3716	)	,
(	3715	)	,
(	3713	)	,
(	3712	)	,
(	3711	)	,
(	3710	)	,
(	3708	)	,
(	3707	)	,
(	3706	)	,
(	3705	)	,
(	3704	)	,
(	3702	)	,
(	3701	)	,
(	3700	)	,
(	3699	)	,
(	3697	)	,
(	3696	)	,
(	3695	)	,
(	3694	)	,
(	3692	)	,
(	3691	)	,
(	3690	)	,
(	3689	)	,
(	3687	)	,
(	3686	)	,
(	3685	)	,
(	3684	)	,
(	3683	)	,
(	3681	)	,
(	3680	)	,
(	3679	)	,
(	3678	)	,
(	3676	)	,
(	3675	)	,
(	3674	)	,
(	3673	)	,
(	3671	)	,
(	3670	)	,
(	3669	)	,
(	3668	)	,
(	3667	)	,
(	3665	)	,
(	3664	)	,
(	3663	)	,
(	3662	)	,
(	3660	)	,
(	3659	)	,
(	3658	)	,
(	3657	)	,
(	3655	)	,
(	3654	)	,
(	3653	)	,
(	3652	)	,
(	3650	)	,
(	3649	)	,
(	3648	)	,
(	3647	)	,
(	3646	)	,
(	3644	)	,
(	3643	)	,
(	3642	)	,
(	3641	)	,
(	3639	)	,
(	3638	)	,
(	3637	)	,
(	3636	)	,
(	3634	)	,
(	3633	)	,
(	3632	)	,
(	3631	)	,
(	3629	)	,
(	3628	)	,
(	3627	)	,
(	3626	)	,
(	3625	)	,
(	3623	)	,
(	3622	)	,
(	3621	)	,
(	3620	)	,
(	3618	)	,
(	3617	)	,
(	3616	)	,
(	3615	)	,
(	3613	)	,
(	3612	)	,
(	3611	)	,
(	3610	)	,
(	3609	)	,
(	3607	)	,
(	3606	)	,
(	3605	)	,
(	3604	)	,
(	3602	)	,
(	3601	)	,
(	3600	)	,
(	3599	)	,
(	3597	)	,
(	3596	)	,
(	3595	)	,
(	3594	)	,
(	3592	)	,
(	3591	)	,
(	3590	)	,
(	3589	)	,
(	3588	)	,
(	3586	)	,
(	3585	)	,
(	3584	)	,
(	3583	)	,
(	3581	)	,
(	3580	)	,
(	3579	)	,
(	3578	)	,
(	3576	)	,
(	3575	)	,
(	3574	)	,
(	3573	)	,
(	3571	)	,
(	3570	)	,
(	3569	)	,
(	3568	)	,
(	3567	)	,
(	3565	)	,
(	3564	)	,
(	3563	)	,
(	3562	)	,
(	3560	)	,
(	3559	)	,
(	3558	)	,
(	3557	)	,
(	3555	)	,
(	3554	)	,
(	3553	)	,
(	3552	)	,
(	3551	)	,
(	3549	)	,
(	3548	)	,
(	3547	)	,
(	3546	)	,
(	3544	)	,
(	3543	)	,
(	3542	)	,
(	3541	)	,
(	3539	)	,
(	3538	)	,
(	3537	)	,
(	3536	)	,
(	3534	)	,
(	3533	)	,
(	3532	)	,
(	3531	)	,
(	3530	)	,
(	3528	)	,
(	3527	)	,
(	3526	)	,
(	3525	)	,
(	3523	)	,
(	3522	)	,
(	3521	)	,
(	3520	)	,
(	3518	)	,
(	3517	)	,
(	3516	)	,
(	3515	)	,
(	3513	)	,
(	3512	)	,
(	3511	)	,
(	3510	)	,
(	3509	)	,
(	3507	)	,
(	3506	)	,
(	3505	)	,
(	3504	)	,
(	3502	)	,
(	3501	)	,
(	3500	)	,
(	3499	)	,
(	3497	)	,
(	3496	)	,
(	3495	)	,
(	3494	)	,
(	3493	)	,
(	3491	)	,
(	3490	)	,
(	3489	)	,
(	3488	)	,
(	3486	)	,
(	3485	)	,
(	3484	)	,
(	3483	)	,
(	3481	)	,
(	3480	)	,
(	3479	)	,
(	3478	)	,
(	3476	)	,
(	3475	)	,
(	3474	)	,
(	3473	)	,
(	3472	)	,
(	3470	)	,
(	3469	)	,
(	3468	)	,
(	3467	)	,
(	3465	)	,
(	3464	)	,
(	3463	)	,
(	3462	)	,
(	3460	)	,
(	3459	)	,
(	3458	)	,
(	3457	)	,
(	3455	)	,
(	3454	)	,
(	3453	)	,
(	3452	)	,
(	3451	)	,
(	3449	)	,
(	3448	)	,
(	3447	)	,
(	3446	)	,
(	3444	)	,
(	3443	)	,
(	3442	)	,
(	3441	)	,
(	3439	)	,
(	3438	)	,
(	3437	)	,
(	3436	)	,
(	3435	)	,
(	3433	)	,
(	3432	)	,
(	3431	)	,
(	3430	)	,
(	3428	)	,
(	3427	)	,
(	3426	)	,
(	3425	)	,
(	3423	)	,
(	3422	)	,
(	3421	)	,
(	3420	)	,
(	3418	)	,
(	3417	)	,
(	3416	)	,
(	3415	)	,
(	3414	)	,
(	3412	)	,
(	3411	)	,
(	3410	)	,
(	3409	)	,
(	3407	)	,
(	3406	)	,
(	3405	)	,
(	3404	)	,
(	3402	)	,
(	3401	)	,
(	3400	)	,
(	3399	)	,
(	3397	)	,
(	3396	)	,
(	3395	)	,
(	3394	)	,
(	3393	)	,
(	3391	)	,
(	3390	)	,
(	3389	)	,
(	3388	)	,
(	3386	)	,
(	3385	)	,
(	3384	)	,
(	3383	)	,
(	3381	)	,
(	3380	)	,
(	3379	)	,
(	3378	)	,
(	3377	)	,
(	3375	)	,
(	3374	)	,
(	3373	)	,
(	3372	)	,
(	3370	)	,
(	3369	)	,
(	3368	)	,
(	3367	)	,
(	3365	)	,
(	3364	)	,
(	3363	)	,
(	3362	)	,
(	3360	)	,
(	3359	)	,
(	3358	)	,
(	3357	)	,
(	3356	)	,
(	3354	)	,
(	3353	)	,
(	3352	)	,
(	3351	)	,
(	3349	)	,
(	3348	)	,
(	3347	)	,
(	3346	)	,
(	3344	)	,
(	3343	)	,
(	3342	)	,
(	3341	)	,
(	3339	)	,
(	3338	)	,
(	3337	)	,
(	3336	)	,
(	3335	)	,
(	3333	)	,
(	3332	)	,
(	3331	)	,
(	3330	)	,
(	3328	)	,
(	3327	)	,
(	3326	)	,
(	3325	)	,
(	3323	)	,
(	3322	)	,
(	3321	)	,
(	3320	)	,
(	3319	)	,
(	3317	)	,
(	3316	)	,
(	3315	)	,
(	3314	)	,
(	3312	)	,
(	3311	)	,
(	3310	)	,
(	3309	)	,
(	3307	)	,
(	3306	)	,
(	3305	)	,
(	3304	)	,
(	3302	)	,
(	3301	)	,
(	3300	)	,
(	3299	)	,
(	3298	)	,
(	3296	)	,
(	3295	)	,
(	3294	)	,
(	3293	)	,
(	3291	)	,
(	3290	)	,
(	3289	)	,
(	3288	)	,
(	3286	)	,
(	3285	)	,
(	3284	)	,
(	3283	)	,
(	3281	)	,
(	3280	)	,
(	3279	)	,
(	3278	)	,
(	3277	)	,
(	3275	)	,
(	3274	)	,
(	3273	)	,
(	3272	)	,
(	3270	)	,
(	3269	)	,
(	3268	)	,
(	3267	)	,
(	3265	)	,
(	3264	)	,
(	3263	)	,
(	3262	)	,
(	3261	)	,
(	3259	)	,
(	3258	)	,
(	3257	)	,
(	3256	)	,
(	3254	)	,
(	3253	)	,
(	3252	)	,
(	3251	)	,
(	3249	)	,
(	3248	)	,
(	3247	)	,
(	3246	)	,
(	3244	)	,
(	3243	)	,
(	3242	)	,
(	3241	)	,
(	3240	)	,
(	3238	)	,
(	3237	)	,
(	3236	)	,
(	3235	)	,
(	3233	)	,
(	3232	)	,
(	3231	)	,
(	3230	)	,
(	3228	)	,
(	3227	)	,
(	3226	)	,
(	3225	)	,
(	3223	)	,
(	3222	)	,
(	3221	)	,
(	3220	)	,
(	3219	)	,
(	3217	)	,
(	3216	)	,
(	3215	)	,
(	3214	)	,
(	3212	)	,
(	3211	)	,
(	3210	)	,
(	3209	)	,
(	3207	)	,
(	3206	)	,
(	3205	)	,
(	3204	)	,
(	3203	)	,
(	3201	)	,
(	3200	)	,
(	3199	)	,
(	3198	)	,
(	3196	)	,
(	3195	)	,
(	3194	)	,
(	3193	)	,
(	3191	)	,
(	3190	)	,
(	3189	)	,
(	3188	)	,
(	3186	)	,
(	3185	)	,
(	3184	)	,
(	3183	)	,
(	3182	)	,
(	3180	)	,
(	3179	)	,
(	3178	)	,
(	3177	)	,
(	3175	)	,
(	3174	)	,
(	3173	)	,
(	3172	)	,
(	3170	)	,
(	3169	)	,
(	3168	)	,
(	3167	)	,
(	3165	)	,
(	3164	)	,
(	3163	)	,
(	3162	)	,
(	3161	)	,
(	3159	)	,
(	3158	)	,
(	3157	)	,
(	3156	)	,
(	3154	)	,
(	3153	)	,
(	3152	)	,
(	3151	)	,
(	3149	)	,
(	3148	)	,
(	3147	)	,
(	3146	)	,
(	3145	)	,
(	3143	)	,
(	3142	)	,
(	3141	)	,
(	3140	)	,
(	3138	)	,
(	3137	)	,
(	3136	)	,
(	3135	)	,
(	3133	)	,
(	3132	)	,
(	3131	)	,
(	3130	)	,
(	3128	)	,
(	3127	)	,
(	3126	)	,
(	3125	)	,
(	3124	)	,
(	3122	)	,
(	3121	)	,
(	3120	)	,
(	3119	)	,
(	3117	)	,
(	3116	)	,
(	3115	)	,
(	3114	)	,
(	3112	)	,
(	3111	)	,
(	3110	)	,
(	3109	)	,
(	3107	)	,
(	3106	)	,
(	3105	)	,
(	3104	)	,
(	3103	)	,
(	3101	)	,
(	3100	)	,
(	3099	)	,
(	3098	)	,
(	3096	)	,
(	3095	)	,
(	3094	)	,
(	3093	)	,
(	3091	)	,
(	3090	)	,
(	3089	)	,
(	3088	)	,
(	3087	)	,
(	3085	)	,
(	3084	)	,
(	3083	)	,
(	3082	)	,
(	3080	)	,
(	3079	)	,
(	3078	)	,
(	3077	)	,
(	3075	)	,
(	3074	)	,
(	3073	)	,
(	3072	)	,
(	3070	)	,
(	3069	)	,
(	3068	)	,
(	3067	)	,
(	3066	)	,
(	3064	)	,
(	3063	)	,
(	3062	)	,
(	3061	)	,
(	3059	)	,
(	3058	)	,
(	3057	)	,
(	3056	)	,
(	3054	)	,
(	3053	)	,
(	3052	)	,
(	3051	)	,
(	3049	)	,
(	3048	)	,
(	3047	)	,
(	3046	)	,
(	3045	)	,
(	3043	)	,
(	3042	)	,
(	3041	)	,
(	3040	)	,
(	3038	)	,
(	3037	)	,
(	3036	)	,
(	3035	)	,
(	3033	)	,
(	3032	)	,
(	3031	)	,
(	3030	)	,
(	3029	)	,
(	3027	)	,
(	3026	)	,
(	3025	)	,
(	3024	)	,
(	3022	)	,
(	3021	)	,
(	3020	)	,
(	3019	)	,
(	3017	)	,
(	3016	)	,
(	3015	)	,
(	3014	)	,
(	3012	)	,
(	3011	)	,
(	3010	)	,
(	3009	)	,
(	3008	)	,
(	3006	)	,
(	3005	)	,
(	3004	)	,
(	3003	)	,
(	3001	)	,
(	3000	)	,
(	2999	)	,
(	2998	)	,
(	2996	)	,
(	2995	)	,
(	2994	)	,
(	2993	)	,
(	2991	)	,
(	2990	)	,
(	2989	)	,
(	2988	)	,
(	2987	)	,
(	2985	)	,
(	2984	)	,
(	2983	)	,
(	2982	)	,
(	2980	)	,
(	2979	)	,
(	2978	)	,
(	2977	)	,
(	2975	)	,
(	2974	)	,
(	2973	)	,
(	2972	)	,
(	2971	)	,
(	2969	)	,
(	2968	)	,
(	2967	)	,
(	2966	)	,
(	2964	)	,
(	2963	)	,
(	2962	)	,
(	2961	)	,
(	2959	)	,
(	2958	)	,
(	2957	)	,
(	2956	)	,
(	2954	)	,
(	2953	)	,
(	2952	)	,
(	2951	)	,
(	2950	)	,
(	2948	)	,
(	2947	)	,
(	2946	)	,
(	2945	)	,
(	2943	)	,
(	2942	)	,
(	2941	)	,
(	2940	)	,
(	2938	)	,
(	2937	)	,
(	2936	)	,
(	2935	)	,
(	2933	)	,
(	2932	)	,
(	2931	)	,
(	2930	)	,
(	2929	)	,
(	2927	)	,
(	2926	)	,
(	2925	)	,
(	2924	)	,
(	2922	)	,
(	2921	)	,
(	2920	)	,
(	2919	)	,
(	2917	)	,
(	2916	)	,
(	2915	)	,
(	2914	)	,
(	2913	)	,
(	2911	)	,
(	2910	)	,
(	2909	)	,
(	2908	)	,
(	2906	)	,
(	2905	)	,
(	2904	)	,
(	2903	)	,
(	2901	)	,
(	2900	)	,
(	2899	)	,
(	2898	)	,
(	2896	)	,
(	2895	)	,
(	2894	)	,
(	2893	)	,
(	2892	)	,
(	2890	)	,
(	2889	)	,
(	2888	)	,
(	2887	)	,
(	2885	)	,
(	2884	)	,
(	2883	)	,
(	2882	)	,
(	2880	)	,
(	2879	)	,
(	2878	)	,
(	2877	)	,
(	2875	)	,
(	2874	)	,
(	2873	)	,
(	2872	)	,
(	2871	)	,
(	2869	)	,
(	2868	)	,
(	2867	)	,
(	2866	)	,
(	2864	)	,
(	2863	)	,
(	2862	)	,
(	2861	)	,
(	2859	)	,
(	2858	)	,
(	2857	)	,
(	2856	)	,
(	2855	)	,
(	2853	)	,
(	2852	)	,
(	2851	)	,
(	2850	)	,
(	2848	)	,
(	2847	)	,
(	2846	)	,
(	2845	)	,
(	2843	)	,
(	2842	)	,
(	2841	)	,
(	2840	)	,
(	2838	)	,
(	2837	)	,
(	2836	)	,
(	2835	)	,
(	2834	)	,
(	2832	)	,
(	2831	)	,
(	2830	)	,
(	2829	)	,
(	2827	)	,
(	2826	)	,
(	2825	)	,
(	2824	)	,
(	2822	)	,
(	2821	)	,
(	2820	)	,
(	2819	)	,
(	2817	)	,
(	2816	)	,
(	2815	)	,
(	2814	)	,
(	2813	)	,
(	2811	)	,
(	2810	)	,
(	2809	)	,
(	2808	)	,
(	2806	)	,
(	2805	)	,
(	2804	)	,
(	2803	)	,
(	2801	)	,
(	2800	)	,
(	2799	)	,
(	2798	)	,
(	2797	)	,
(	2795	)	,
(	2794	)	,
(	2793	)	,
(	2792	)	,
(	2790	)	,
(	2789	)	,
(	2788	)	,
(	2787	)	,
(	2785	)	,
(	2784	)	,
(	2783	)	,
(	2782	)	,
(	2780	)	,
(	2779	)	,
(	2778	)	,
(	2777	)	,
(	2776	)	,
(	2774	)	,
(	2773	)	,
(	2772	)	,
(	2771	)	,
(	2769	)	,
(	2768	)	,
(	2767	)	,
(	2766	)	,
(	2764	)	,
(	2763	)	,
(	2762	)	,
(	2761	)	,
(	2759	)	,
(	2758	)	,
(	2757	)	,
(	2756	)	,
(	2755	)	,
(	2753	)	,
(	2752	)	,
(	2751	)	,
(	2750	)	,
(	2748	)	,
(	2747	)	,
(	2746	)	,
(	2745	)	,
(	2743	)	,
(	2742	)	,
(	2741	)	,
(	2740	)	,
(	2739	)	,
(	2737	)	,
(	2736	)	,
(	2735	)	,
(	2734	)	,
(	2732	)	,
(	2731	)	,
(	2730	)	,
(	2729	)	,
(	2727	)	,
(	2726	)	,
(	2725	)	,
(	2724	)	,
(	2722	)	,
(	2721	)	,
(	2720	)	,
(	2719	)	,
(	2718	)	,
(	2716	)	,
(	2715	)	,
(	2714	)	,
(	2713	)	,
(	2711	)	,
(	2710	)	,
(	2709	)	,
(	2708	)	,
(	2706	)	,
(	2705	)	,
(	2704	)	,
(	2703	)	,
(	2701	)	,
(	2700	)	,
(	2699	)	,
(	2698	)	,
(	2697	)	,
(	2695	)	,
(	2694	)	,
(	2693	)	,
(	2692	)	,
(	2690	)	,
(	2689	)	,
(	2688	)	,
(	2687	)	,
(	2685	)	,
(	2684	)	,
(	2683	)	,
(	2682	)	,
(	2681	)	,
(	2679	)	,
(	2678	)	,
(	2677	)	,
(	2676	)	,
(	2674	)	,
(	2673	)	,
(	2672	)	,
(	2671	)	,
(	2669	)	,
(	2668	)	,
(	2667	)	,
(	2666	)	,
(	2664	)	,
(	2663	)	,
(	2662	)	,
(	2661	)	,
(	2660	)	,
(	2658	)	,
(	2657	)	,
(	2656	)	,
(	2655	)	,
(	2653	)	,
(	2652	)	,
(	2651	)	,
(	2650	)	,
(	2648	)	,
(	2647	)	,
(	2646	)	,
(	2645	)	,
(	2643	)	,
(	2642	)	,
(	2641	)	,
(	2640	)	,
(	2639	)	,
(	2637	)	,
(	2636	)	,
(	2635	)	,
(	2634	)	,
(	2632	)	,
(	2631	)	,
(	2630	)	,
(	2629	)	,
(	2627	)	,
(	2626	)	,
(	2625	)	,
(	2624	)	,
(	2623	)	,
(	2621	)	,
(	2620	)	,
(	2619	)	,
(	2618	)	,
(	2616	)	,
(	2615	)	,
(	2614	)	,
(	2613	)	,
(	2611	)	,
(	2610	)	,
(	2609	)	,
(	2608	)	,
(	2606	)	,
(	2605	)	,
(	2604	)	,
(	2603	)	,
(	2602	)	,
(	2600	)	,
(	2599	)	,
(	2598	)	,
(	2597	)	,
(	2595	)	,
(	2594	)	,
(	2593	)	,
(	2592	)	,
(	2590	)	,
(	2589	)	,
(	2588	)	,
(	2587	)	,
(	2585	)	,
(	2584	)	,
(	2583	)	,
(	2582	)	,
(	2581	)	,
(	2579	)	,
(	2578	)	,
(	2577	)	,
(	2576	)	,
(	2574	)	,
(	2573	)	,
(	2572	)	,
(	2571	)	,
(	2569	)	,
(	2568	)	,
(	2567	)	,
(	2566	)	,
(	2565	)	,
(	2563	)	,
(	2562	)	,
(	2561	)	,
(	2560	)	,
(	2558	)	,
(	2557	)	,
(	2556	)	,
(	2555	)	,
(	2553	)	,
(	2552	)	,
(	2551	)	,
(	2550	)	,
(	2548	)	,
(	2547	)	,
(	2546	)	,
(	2545	)	,
(	2544	)	,
(	2542	)	,
(	2541	)	,
(	2540	)	,
(	2539	)	,
(	2537	)	,
(	2536	)	,
(	2535	)	,
(	2534	)	,
(	2532	)	,
(	2531	)	,
(	2530	)	,
(	2529	)	,
(	2527	)	,
(	2526	)	,
(	2525	)	,
(	2524	)	,
(	2523	)	,
(	2521	)	,
(	2520	)	,
(	2519	)	,
(	2518	)	,
(	2516	)	,
(	2515	)	,
(	2514	)	,
(	2513	)	,
(	2511	)	,
(	2510	)	,
(	2509	)	,
(	2508	)	,
(	2507	)	,
(	2505	)	,
(	2504	)	,
(	2503	)	,
(	2502	)	,
(	2500	)	,
(	2499	)	,
(	2498	)	,
(	2497	)	,
(	2495	)	,
(	2494	)	,
(	2493	)	,
(	2492	)	,
(	2490	)	,
(	2489	)	,
(	2488	)	,
(	2487	)	,
(	2486	)	,
(	2484	)	,
(	2483	)	,
(	2482	)	,
(	2481	)	,
(	2479	)	,
(	2478	)	,
(	2477	)	,
(	2476	)	,
(	2474	)	,
(	2473	)	,
(	2472	)	,
(	2471	)	,
(	2469	)	,
(	2468	)	,
(	2467	)	,
(	2466	)	,
(	2465	)	,
(	2463	)	,
(	2462	)	,
(	2461	)	,
(	2460	)	,
(	2458	)	,
(	2457	)	,
(	2456	)	,
(	2455	)	,
(	2453	)	,
(	2452	)	,
(	2451	)	,
(	2450	)	,
(	2449	)	,
(	2447	)	,
(	2446	)	,
(	2445	)	,
(	2444	)	,
(	2442	)	,
(	2441	)	,
(	2440	)	,
(	2439	)	,
(	2437	)	,
(	2436	)	,
(	2435	)	,
(	2434	)	,
(	2432	)	,
(	2431	)	,
(	2430	)	,
(	2429	)	,
(	2428	)	,
(	2426	)	,
(	2425	)	,
(	2424	)	,
(	2423	)	,
(	2421	)	,
(	2420	)	,
(	2419	)	,
(	2418	)	,
(	2416	)	,
(	2415	)	,
(	2414	)	,
(	2413	)	,
(	2411	)	,
(	2410	)	,
(	2409	)	,
(	2408	)	,
(	2407	)	,
(	2405	)	,
(	2404	)	,
(	2403	)	,
(	2402	)	,
(	2400	)	,
(	2399	)	,
(	2398	)	,
(	2397	)	,
(	2395	)	,
(	2394	)	,
(	2393	)	,
(	2392	)	,
(	2391	)	,
(	2389	)	,
(	2388	)	,
(	2387	)	,
(	2386	)	,
(	2384	)	,
(	2383	)	,
(	2382	)	,
(	2381	)	,
(	2379	)	,
(	2378	)	,
(	2377	)	,
(	2376	)	,
(	2374	)	,
(	2373	)	,
(	2372	)	,
(	2371	)	,
(	2370	)	,
(	2368	)	,
(	2367	)	,
(	2366	)	,
(	2365	)	,
(	2363	)	,
(	2362	)	,
(	2361	)	,
(	2360	)	,
(	2358	)	,
(	2357	)	,
(	2356	)	,
(	2355	)	,
(	2353	)	,
(	2352	)	,
(	2351	)	,
(	2350	)	,
(	2349	)	,
(	2347	)	,
(	2346	)	,
(	2345	)	,
(	2344	)	,
(	2342	)	,
(	2341	)	,
(	2340	)	,
(	2339	)	,
(	2337	)	,
(	2336	)	,
(	2335	)	,
(	2334	)	,
(	2333	)	,
(	2331	)	,
(	2330	)	,
(	2329	)	,
(	2328	)	,
(	2326	)	,
(	2325	)	,
(	2324	)	,
(	2323	)	,
(	2321	)	,
(	2320	)	,
(	2319	)	,
(	2318	)	,
(	2316	)	,
(	2315	)	,
(	2314	)	,
(	2313	)	,
(	2312	)	,
(	2310	)	,
(	2309	)	,
(	2308	)	,
(	2307	)	,
(	2305	)	,
(	2304	)	,
(	2303	)	,
(	2302	)	,
(	2300	)	,
(	2299	)	,
(	2298	)	,
(	2297	)	,
(	2295	)	,
(	2294	)	,
(	2293	)	,
(	2292	)	,
(	2291	)	,
(	2289	)	,
(	2288	)	,
(	2287	)	,
(	2286	)	,
(	2284	)	,
(	2283	)	,
(	2282	)	,
(	2281	)	,
(	2279	)	,
(	2278	)	,
(	2277	)	,
(	2276	)	,
(	2275	)	,
(	2273	)	,
(	2272	)	,
(	2271	)	,
(	2270	)	,
(	2268	)	,
(	2267	)	,
(	2266	)	,
(	2265	)	,
(	2263	)	,
(	2262	)	,
(	2261	)	,
(	2260	)	,
(	2258	)	,
(	2257	)	,
(	2256	)	,
(	2255	)	,
(	2254	)	,
(	2252	)	,
(	2251	)	,
(	2250	)	,
(	2249	)	,
(	2247	)	,
(	2246	)	,
(	2245	)	,
(	2244	)	,
(	2242	)	,
(	2241	)	,
(	2240	)	,
(	2239	)	,
(	2237	)	,
(	2236	)	,
(	2235	)	,
(	2234	)	,
(	2233	)	,
(	2231	)	,
(	2230	)	,
(	2229	)	,
(	2228	)	,
(	2226	)	,
(	2225	)	,
(	2224	)	,
(	2223	)	,
(	2221	)	,
(	2220	)	,
(	2219	)	,
(	2218	)	,
(	2217	)	,
(	2215	)	,
(	2214	)	,
(	2213	)	,
(	2212	)	,
(	2210	)	,
(	2209	)	,
(	2208	)	,
(	2207	)	,
(	2205	)	,
(	2204	)	,
(	2203	)	,
(	2202	)	,
(	2200	)	,
(	2199	)	,
(	2198	)	,
(	2197	)	,
(	2196	)	,
(	2194	)	,
(	2193	)	,
(	2192	)	,
(	2191	)	,
(	2189	)	,
(	2188	)	,
(	2187	)	,
(	2186	)	,
(	2184	)	,
(	2183	)	,
(	2182	)	,
(	2181	)	,
(	2179	)	,
(	2178	)	,
(	2177	)	,
(	2176	)	,
(	2175	)	,
(	2173	)	,
(	2172	)	,
(	2171	)	,
(	2170	)	,
(	2168	)	,
(	2167	)	,
(	2166	)	,
(	2165	)	,
(	2163	)	,
(	2162	)	,
(	2161	)	,
(	2160	)	,
(	2159	)	,
(	2157	)	,
(	2156	)	,
(	2155	)	,
(	2154	)	,
(	2152	)	,
(	2151	)	,
(	2150	)	,
(	2149	)	,
(	2147	)	,
(	2146	)	,
(	2145	)	,
(	2144	)	,
(	2142	)	,
(	2141	)	,
(	2140	)	,
(	2139	)	,
(	2138	)	,
(	2136	)	,
(	2135	)	,
(	2134	)	,
(	2133	)	,
(	2131	)	,
(	2130	)	,
(	2129	)	,
(	2128	)	,
(	2126	)	,
(	2125	)	,
(	2124	)	,
(	2123	)	,
(	2121	)	,
(	2120	)	,
(	2119	)	,
(	2118	)	,
(	2117	)	,
(	2115	)	,
(	2114	)	,
(	2113	)	,
(	2112	)	,
(	2110	)	,
(	2109	)	,
(	2108	)	,
(	2107	)	,
(	2105	)	,
(	2104	)	,
(	2103	)	,
(	2102	)	,
(	2101	)	,
(	2099	)	,
(	2098	)	,
(	2097	)	,
(	2096	)	,
(	2094	)	,
(	2093	)	,
(	2092	)	,
(	2091	)	,
(	2089	)	,
(	2088	)	,
(	2087	)	,
(	2086	)	,
(	2084	)	,
(	2083	)	,
(	2082	)	,
(	2081	)	,
(	2080	)	,
(	2078	)	,
(	2077	)	,
(	2076	)	,
(	2075	)	,
(	2073	)	,
(	2072	)	,
(	2071	)	,
(	2070	)	,
(	2068	)	,
(	2067	)	,
(	2066	)	,
(	2065	)	,
(	2063	)	,
(	2062	)	,
(	2061	)	,
(	2060	)	,
(	2059	)	,
(	2057	)	,
(	2056	)	,
(	2055	)	,
(	2054	)	,
(	2052	)	,
(	2051	)	,
(	2050	)	,
(	2049	)	,
(	2047	)	,
(	2046	)	,
(	2045	)	,
(	2044	)	,
(	2043	)	,
(	2041	)	,
(	2040	)	,
(	2039	)	,
(	2038	)	,
(	2036	)	,
(	2035	)	,
(	2034	)	,
(	2033	)	,
(	2031	)	,
(	2030	)	,
(	2029	)	,
(	2028	)	,
(	2026	)	,
(	2025	)	,
(	2024	)	,
(	2023	)	,
(	2022	)	,
(	2020	)	,
(	2019	)	,
(	2018	)	,
(	2017	)	,
(	2015	)	,
(	2014	)	,
(	2013	)	,
(	2012	)	,
(	2010	)	,
(	2009	)	,
(	2008	)	,
(	2007	)	,
(	2005	)	,
(	2004	)	,
(	2003	)	,
(	2002	)	,
(	2001	)	,
(	1999	)	,
(	1998	)	,
(	1997	)	,
(	1996	)	,
(	1994	)	,
(	1993	)	,
(	1992	)	,
(	1991	)	,
(	1989	)	,
(	1988	)	,
(	1987	)	,
(	1986	)	,
(	1985	)	,
(	1983	)	,
(	1982	)	,
(	1981	)	,
(	1980	)	,
(	1978	)	,
(	1977	)	,
(	1976	)	,
(	1975	)	,
(	1973	)	,
(	1972	)	,
(	1971	)	,
(	1970	)	,
(	1968	)	,
(	1967	)	,
(	1966	)	,
(	1965	)	,
(	1964	)	,
(	1962	)	,
(	1961	)	,
(	1960	)	,
(	1959	)	,
(	1957	)	,
(	1956	)	,
(	1955	)	,
(	1954	)	,
(	1952	)	,
(	1951	)	,
(	1950	)	,
(	1949	)	,
(	1947	)	,
(	1946	)	,
(	1945	)	,
(	1944	)	,
(	1943	)	,
(	1941	)	,
(	1940	)	,
(	1939	)	,
(	1938	)	,
(	1936	)	,
(	1935	)	,
(	1934	)	,
(	1933	)	,
(	1931	)	,
(	1930	)	,
(	1929	)	,
(	1928	)	,
(	1927	)	,
(	1925	)	,
(	1924	)	,
(	1923	)	,
(	1922	)	,
(	1920	)	,
(	1919	)	,
(	1918	)	,
(	1917	)	,
(	1915	)	,
(	1914	)	,
(	1913	)	,
(	1912	)	,
(	1910	)	,
(	1909	)	,
(	1908	)	,
(	1907	)	,
(	1906	)	,
(	1904	)	,
(	1903	)	,
(	1902	)	,
(	1901	)	,
(	1899	)	,
(	1898	)	,
(	1897	)	,
(	1896	)	,
(	1894	)	,
(	1893	)	,
(	1892	)	,
(	1891	)	,
(	1889	)	,
(	1888	)	,
(	1887	)	,
(	1886	)	,
(	1885	)	,
(	1883	)	,
(	1882	)	,
(	1881	)	,
(	1880	)	,
(	1878	)	,
(	1877	)	,
(	1876	)	,
(	1875	)	,
(	1873	)	,
(	1872	)	,
(	1871	)	,
(	1870	)	,
(	1869	)	,
(	1867	)	,
(	1866	)	,
(	1865	)	,
(	1864	)	,
(	1862	)	,
(	1861	)	,
(	1860	)	,
(	1859	)	,
(	1857	)	,
(	1856	)	,
(	1855	)	,
(	1854	)	,
(	1852	)	,
(	1851	)	,
(	1850	)	,
(	1849	)	,
(	1848	)	,
(	1846	)	,
(	1845	)	,
(	1844	)	,
(	1843	)	,
(	1841	)	,
(	1840	)	,
(	1839	)	,
(	1838	)	,
(	1836	)	,
(	1835	)	,
(	1834	)	,
(	1833	)	,
(	1831	)	,
(	1830	)	,
(	1829	)	,
(	1828	)	,
(	1827	)	,
(	1825	)	,
(	1824	)	,
(	1823	)	,
(	1822	)	,
(	1820	)	,
(	1819	)	,
(	1818	)	,
(	1817	)	,
(	1815	)	,
(	1814	)	,
(	1813	)	,
(	1812	)	,
(	1811	)	,
(	1809	)	,
(	1808	)	,
(	1807	)	,
(	1806	)	,
(	1804	)	,
(	1803	)	,
(	1802	)	,
(	1801	)	,
(	1799	)	,
(	1798	)	,
(	1797	)	,
(	1796	)	,
(	1794	)	,
(	1793	)	,
(	1792	)	,
(	1791	)	,
(	1790	)	,
(	1788	)	,
(	1787	)	,
(	1786	)	,
(	1785	)	,
(	1783	)	,
(	1782	)	,
(	1781	)	,
(	1780	)	,
(	1778	)	,
(	1777	)	,
(	1776	)	,
(	1775	)	,
(	1773	)	,
(	1772	)	,
(	1771	)	,
(	1770	)	,
(	1769	)	,
(	1767	)	,
(	1766	)	,
(	1765	)	,
(	1764	)	,
(	1762	)	,
(	1761	)	,
(	1760	)	,
(	1759	)	,
(	1757	)	,
(	1756	)	,
(	1755	)	,
(	1754	)	,
(	1753	)	,
(	1751	)	,
(	1750	)	,
(	1749	)	,
(	1748	)	,
(	1746	)	,
(	1745	)	,
(	1744	)	,
(	1743	)	,
(	1741	)	,
(	1740	)	,
(	1739	)	,
(	1738	)	,
(	1736	)	,
(	1735	)	,
(	1734	)	,
(	1733	)	,
(	1732	)	,
(	1730	)	,
(	1729	)	,
(	1728	)	,
(	1727	)	,
(	1725	)	,
(	1724	)	,
(	1723	)	,
(	1722	)	,
(	1720	)	,
(	1719	)	,
(	1718	)	,
(	1717	)	,
(	1715	)	,
(	1714	)	,
(	1713	)	,
(	1712	)	,
(	1711	)	,
(	1709	)	,
(	1708	)	,
(	1707	)	,
(	1706	)	,
(	1704	)	,
(	1703	)	,
(	1702	)	,
(	1701	)	,
(	1699	)	,
(	1698	)	,
(	1697	)	,
(	1696	)	,
(	1695	)	,
(	1693	)	,
(	1692	)	,
(	1691	)	,
(	1690	)	,
(	1688	)	,
(	1687	)	,
(	1686	)	,
(	1685	)	,
(	1683	)	,
(	1682	)	,
(	1681	)	,
(	1680	)	,
(	1678	)	,
(	1677	)	,
(	1676	)	,
(	1675	)	,
(	1674	)	,
(	1672	)	,
(	1671	)	,
(	1670	)	,
(	1669	)	,
(	1667	)	,
(	1666	)	,
(	1665	)	,
(	1664	)	,
(	1662	)	,
(	1661	)	,
(	1660	)	,
(	1659	)	,
(	1657	)	,
(	1656	)	,
(	1655	)	,
(	1654	)	,
(	1653	)	,
(	1651	)	,
(	1650	)	,
(	1649	)	,
(	1648	)	,
(	1646	)	,
(	1645	)	,
(	1644	)	,
(	1643	)	,
(	1641	)	,
(	1640	)	,
(	1639	)	,
(	1638	)	,
(	1637	)	,
(	1635	)	,
(	1634	)	,
(	1633	)	,
(	1632	)	,
(	1630	)	,
(	1629	)	,
(	1628	)	,
(	1627	)	,
(	1625	)	,
(	1624	)	,
(	1623	)	,
(	1622	)	,
(	1620	)	,
(	1619	)	,
(	1618	)	,
(	1617	)	,
(	1616	)	,
(	1614	)	,
(	1613	)	,
(	1612	)	,
(	1611	)	,
(	1609	)	,
(	1608	)	,
(	1607	)	,
(	1606	)	,
(	1604	)	,
(	1603	)	,
(	1602	)	,
(	1601	)	,
(	1599	)	,
(	1598	)	,
(	1597	)	,
(	1596	)	,
(	1595	)	,
(	1593	)	,
(	1592	)	,
(	1591	)	,
(	1590	)	,
(	1588	)	,
(	1587	)	,
(	1586	)	,
(	1585	)	,
(	1583	)	,
(	1582	)	,
(	1581	)	,
(	1580	)	,
(	1579	)	,
(	1577	)	,
(	1576	)	,
(	1575	)	,
(	1574	)	,
(	1572	)	,
(	1571	)	,
(	1570	)	,
(	1569	)	,
(	1567	)	,
(	1566	)	,
(	1565	)	,
(	1564	)	,
(	1562	)	,
(	1561	)	,
(	1560	)	,
(	1559	)	,
(	1558	)	,
(	1556	)	,
(	1555	)	,
(	1554	)	,
(	1553	)	,
(	1551	)	,
(	1550	)	,
(	1549	)	,
(	1548	)	,
(	1546	)	,
(	1545	)	,
(	1544	)	,
(	1543	)	,
(	1541	)	,
(	1540	)	,
(	1539	)	,
(	1538	)	,
(	1537	)	,
(	1535	)	,
(	1534	)	,
(	1533	)	,
(	1532	)	,
(	1530	)	,
(	1529	)	,
(	1528	)	,
(	1527	)	,
(	1525	)	,
(	1524	)	,
(	1523	)	,
(	1522	)	,
(	1521	)	,
(	1519	)	,
(	1518	)	,
(	1517	)	,
(	1516	)	,
(	1514	)	,
(	1513	)	,
(	1512	)	,
(	1511	)	,
(	1509	)	,
(	1508	)	,
(	1507	)	,
(	1506	)	,
(	1504	)	,
(	1503	)	,
(	1502	)	,
(	1501	)	,
(	1500	)	,
(	1498	)	,
(	1497	)	,
(	1496	)	,
(	1495	)	,
(	1493	)	,
(	1492	)	,
(	1491	)	,
(	1490	)	,
(	1488	)	,
(	1487	)	,
(	1486	)	,
(	1485	)	,
(	1483	)	,
(	1482	)	,
(	1481	)	,
(	1480	)	,
(	1479	)	,
(	1477	)	,
(	1476	)	,
(	1475	)	,
(	1474	)	,
(	1472	)	,
(	1471	)	,
(	1470	)	,
(	1469	)	,
(	1467	)	,
(	1466	)	,
(	1465	)	,
(	1464	)	,
(	1463	)	,
(	1461	)	,
(	1460	)	,
(	1459	)	,
(	1458	)	,
(	1456	)	,
(	1455	)	,
(	1454	)	,
(	1453	)	,
(	1451	)	,
(	1450	)	,
(	1449	)	,
(	1448	)	,
(	1446	)	,
(	1445	)	,
(	1444	)	,
(	1443	)	,
(	1442	)	,
(	1440	)	,
(	1439	)	,
(	1438	)	,
(	1437	)	,
(	1435	)	,
(	1434	)	,
(	1433	)	,
(	1432	)	,
(	1430	)	,
(	1429	)	,
(	1428	)	,
(	1427	)	,
(	1425	)	,
(	1424	)	,
(	1423	)	,
(	1422	)	,
(	1421	)	,
(	1419	)	,
(	1418	)	,
(	1417	)	,
(	1416	)	,
(	1414	)	,
(	1413	)	,
(	1412	)	,
(	1411	)	,
(	1409	)	,
(	1408	)	,
(	1407	)	,
(	1406	)	,
(	1405	)	,
(	1403	)	,
(	1402	)	,
(	1401	)	,
(	1400	)	,
(	1398	)	,
(	1397	)	,
(	1396	)	,
(	1395	)	,
(	1393	)	,
(	1392	)	,
(	1391	)	,
(	1390	)	,
(	1388	)	,
(	1387	)	,
(	1386	)	,
(	1385	)	,
(	1384	)	,
(	1382	)	,
(	1381	)	,
(	1380	)	,
(	1379	)	,
(	1377	)	,
(	1376	)	,
(	1375	)	,
(	1374	)	,
(	1372	)	,
(	1371	)	,
(	1370	)	,
(	1369	)	,
(	1367	)	,
(	1366	)	,
(	1365	)	,
(	1364	)	,
(	1363	)	,
(	1361	)	,
(	1360	)	,
(	1359	)	,
(	1358	)	,
(	1356	)	,
(	1355	)	,
(	1354	)	,
(	1353	)	,
(	1351	)	,
(	1350	)	,
(	1349	)	,
(	1348	)	,
(	1347	)	,
(	1345	)	,
(	1344	)	,
(	1343	)	,
(	1342	)	,
(	1340	)	,
(	1339	)	,
(	1338	)	,
(	1337	)	,
(	1335	)	,
(	1334	)	,
(	1333	)	,
(	1332	)	,
(	1330	)	,
(	1329	)	,
(	1328	)	,
(	1327	)	,
(	1326	)	,
(	1324	)	,
(	1323	)	,
(	1322	)	,
(	1321	)	,
(	1319	)	,
(	1318	)	,
(	1317	)	,
(	1316	)	,
(	1314	)	,
(	1313	)	,
(	1312	)	,
(	1311	)	,
(	1309	)	,
(	1308	)	,
(	1307	)	,
(	1306	)	,
(	1305	)	,
(	1303	)	,
(	1302	)	,
(	1301	)	,
(	1300	)	,
(	1298	)	,
(	1297	)	,
(	1296	)	,
(	1295	)	,
(	1293	)	,
(	1292	)	,
(	1291	)	,
(	1290	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1285	)	,
(	1284	)	,
(	1282	)	,
(	1281	)	,
(	1280	)	,
(	1279	)	,
(	1277	)	,
(	1276	)	,
(	1275	)	,
(	1274	)	,
(	1272	)	,
(	1271	)	,
(	1270	)	,
(	1269	)	,
(	1268	)	,
(	1266	)	,
(	1265	)	,
(	1264	)	,
(	1263	)	,
(	1261	)	,
(	1260	)	,
(	1259	)	,
(	1258	)	,
(	1256	)	,
(	1255	)	,
(	1254	)	,
(	1253	)	,
(	1251	)	,
(	1250	)	,
(	1249	)	,
(	1248	)	,
(	1247	)	,
(	1245	)	,
(	1244	)	,
(	1243	)	,
(	1242	)	,
(	1240	)	,
(	1239	)	,
(	1238	)	,
(	1237	)	,
(	1235	)	,
(	1234	)	,
(	1233	)	,
(	1232	)	,
(	1231	)	,
(	1229	)	,
(	1228	)	,
(	1227	)	,
(	1226	)	,
(	1224	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1217	)	,
(	1216	)	,
(	1214	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1210	)	,
(	1208	)	,
(	1207	)	,
(	1206	)	,
(	1205	)	,
(	1203	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1196	)	,
(	1195	)	,
(	1193	)	,
(	1192	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1184	)	,
(	1182	)	,
(	1181	)	,
(	1180	)	,
(	1179	)	,
(	1177	)	,
(	1176	)	,
(	1175	)	,
(	1174	)	,
(	1173	)	,
(	1171	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1152	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1135	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1129	)	,
(	1128	)	,
(	1127	)	,
(	1126	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1121	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1113	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1103	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1089	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	994	)	,
(	992	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	982	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	976	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	968	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	963	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	952	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	947	)	,
(	945	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	941	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	936	)	,
(	934	)	,
(	933	)	,
(	932	)	,
(	931	)	,
(	929	)	,
(	928	)	,
(	927	)	,
(	926	)	,
(	924	)	,
(	923	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	918	)	,
(	917	)	,
(	916	)	,
(	915	)	,
(	913	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	905	)	,
(	903	)	,
(	902	)	,
(	901	)	,
(	900	)	,
(	899	)	,
(	897	)	,
(	896	)	,
(	895	)	,
(	894	)	,
(	892	)	,
(	891	)	,
(	890	)	,
(	889	)	,
(	887	)	,
(	886	)	,
(	885	)	,
(	884	)	,
(	883	)	,
(	881	)	,
(	880	)	,
(	879	)	,
(	878	)	,
(	876	)	,
(	875	)	,
(	874	)	,
(	873	)	,
(	871	)	,
(	870	)	,
(	869	)	,
(	868	)	,
(	866	)	,
(	865	)	,
(	864	)	,
(	863	)	,
(	862	)	,
(	860	)	,
(	859	)	,
(	858	)	,
(	857	)	,
(	855	)	,
(	854	)	,
(	853	)	,
(	852	)	,
(	850	)	,
(	849	)	,
(	848	)	,
(	847	)	,
(	845	)	,
(	844	)	,
(	843	)	,
(	842	)	,
(	841	)	,
(	839	)	,
(	838	)	,
(	837	)	,
(	836	)	,
(	834	)	,
(	833	)	,
(	832	)	,
(	831	)	,
(	829	)	,
(	828	)	,
(	827	)	,
(	826	)	,
(	825	)	,
(	823	)	,
(	822	)	,
(	821	)	,
(	820	)	,
(	818	)	,
(	817	)	,
(	816	)	,
(	815	)	,
(	813	)	,
(	812	)	,
(	811	)	,
(	810	)	,
(	808	)	,
(	807	)	,
(	806	)	,
(	805	)	,
(	804	)	,
(	802	)	,
(	801	)	,
(	800	)	,
(	799	)	,
(	797	)	,
(	796	)	,
(	795	)	,
(	794	)	,
(	792	)	,
(	791	)	,
(	790	)	,
(	789	)	,
(	787	)	,
(	786	)	,
(	785	)	,
(	784	)	,
(	783	)	,
(	781	)	,
(	780	)	,
(	779	)	,
(	778	)	,
(	776	)	,
(	775	)	,
(	774	)	,
(	773	)	,
(	771	)	,
(	770	)	,
(	769	)	,
(	768	)	,
(	767	)	,
(	765	)	,
(	764	)	,
(	763	)	,
(	762	)	,
(	760	)	,
(	759	)	,
(	758	)	,
(	757	)	,
(	755	)	,
(	754	)	,
(	753	)	,
(	752	)	,
(	750	)	,
(	749	)	,
(	748	)	,
(	747	)	,
(	746	)	,
(	744	)	,
(	743	)	,
(	742	)	,
(	741	)	,
(	739	)	,
(	738	)	,
(	737	)	,
(	736	)	,
(	734	)	,
(	733	)	,
(	732	)	,
(	731	)	,
(	729	)	,
(	728	)	,
(	727	)	,
(	726	)	,
(	725	)	,
(	723	)	,
(	722	)	,
(	721	)	,
(	720	)	,
(	718	)	,
(	717	)	,
(	716	)	,
(	715	)	,
(	713	)	,
(	712	)	,
(	711	)	,
(	710	)	,
(	709	)	,
(	707	)	,
(	706	)	,
(	705	)	,
(	704	)	,
(	702	)	,
(	701	)	,
(	700	)	,
(	699	)	,
(	697	)	,
(	696	)	,
(	695	)	,
(	694	)	,
(	692	)	,
(	691	)	,
(	690	)	,
(	689	)	,
(	688	)	,
(	686	)	,
(	685	)	,
(	684	)	,
(	683	)	,
(	681	)	,
(	680	)	,
(	679	)	,
(	678	)	,
(	676	)	,
(	675	)	,
(	674	)	,
(	673	)	,
(	671	)	,
(	670	)	,
(	669	)	,
(	668	)	,
(	667	)	,
(	665	)	,
(	664	)	,
(	663	)	,
(	662	)	,
(	660	)	,
(	659	)	,
(	658	)	,
(	657	)	,
(	655	)	,
(	654	)	,
(	653	)	,
(	652	)	,
(	651	)	,
(	649	)	,
(	648	)	,
(	647	)	,
(	646	)	,
(	644	)	,
(	643	)	,
(	642	)	,
(	641	)	,
(	639	)	,
(	638	)	,
(	637	)	,
(	636	)	,
(	634	)	,
(	633	)	,
(	632	)	,
(	631	)	,
(	630	)	,
(	628	)	,
(	627	)	,
(	626	)	,
(	625	)	,
(	623	)	,
(	622	)	,
(	621	)	,
(	620	)	,
(	618	)	,
(	617	)	,
(	616	)	,
(	615	)	,
(	613	)	,
(	612	)	,
(	611	)	,
(	610	)	,
(	609	)	,
(	607	)	,
(	606	)	,
(	605	)	,
(	604	)	,
(	602	)	,
(	601	)	,
(	600	)	,
(	599	)	,
(	597	)	,
(	596	)	,
(	595	)	,
(	594	)	,
(	593	)	,
(	591	)	,
(	590	)	,
(	589	)	,
(	588	)	,
(	586	)	,
(	585	)	,
(	584	)	,
(	583	)	,
(	581	)	,
(	580	)	,
(	579	)	,
(	578	)	,
(	576	)	,
(	575	)	,
(	574	)	,
(	573	)	,
(	572	)	,
(	570	)	,
(	569	)	,
(	568	)	,
(	567	)	,
(	565	)	,
(	564	)	,
(	563	)	,
(	562	)	,
(	560	)	,
(	559	)	,
(	558	)	,
(	557	)	,
(	555	)	,
(	554	)	,
(	553	)	,
(	552	)	,
(	551	)	,
(	549	)	,
(	548	)	,
(	547	)	,
(	546	)	,
(	544	)	,
(	543	)	,
(	542	)	,
(	541	)	,
(	539	)	,
(	538	)	,
(	537	)	,
(	536	)	,
(	535	)	,
(	533	)	,
(	532	)	,
(	531	)	,
(	530	)	,
(	528	)	,
(	527	)	,
(	526	)	,
(	525	)	,
(	523	)	,
(	522	)	,
(	521	)	,
(	520	)	,
(	518	)	,
(	517	)	,
(	516	)	,
(	515	)	,
(	514	)	,
(	512	)	,
(	511	)	,
(	510	)	,
(	509	)	,
(	507	)	,
(	506	)	,
(	505	)	,
(	504	)	,
(	502	)	,
(	501	)	,
(	500	)	,
(	499	)	,
(	497	)	,
(	496	)	,
(	495	)	,
(	494	)	,
(	493	)	,
(	491	)	,
(	490	)	,
(	489	)	,
(	488	)	,
(	486	)	,
(	485	)	,
(	484	)	,
(	483	)	,
(	481	)	,
(	480	)	,
(	479	)	,
(	478	)	,
(	477	)	,
(	475	)	,
(	474	)	,
(	473	)	,
(	472	)	,
(	470	)	,
(	469	)	,
(	468	)	,
(	467	)	,
(	465	)	,
(	464	)	,
(	463	)	,
(	462	)	,
(	460	)	,
(	459	)	,
(	458	)	,
(	457	)	,
(	456	)	,
(	454	)	,
(	453	)	,
(	452	)	,
(	451	)	,
(	449	)	,
(	448	)	,
(	447	)	,
(	446	)	,
(	444	)	,
(	443	)	,
(	442	)	,
(	441	)	,
(	439	)	,
(	438	)	,
(	437	)	,
(	436	)	,
(	435	)	,
(	433	)	,
(	432	)	,
(	431	)	,
(	430	)	,
(	428	)	,
(	427	)	,
(	426	)	,
(	425	)	,
(	423	)	,
(	422	)	,
(	421	)	,
(	420	)	,
(	419	)	,
(	417	)	,
(	416	)	,
(	415	)	,
(	414	)	,
(	412	)	,
(	411	)	,
(	410	)	,
(	409	)	,
(	407	)	,
(	406	)	,
(	405	)	,
(	404	)	,
(	402	)	,
(	401	)	,
(	400	)	,
(	399	)	,
(	398	)	,
(	396	)	,
(	395	)	,
(	394	)	,
(	393	)	,
(	391	)	,
(	390	)	,
(	389	)	,
(	388	)	,
(	386	)	,
(	385	)	,
(	384	)	,
(	383	)	,
(	381	)	,
(	380	)	,
(	379	)	,
(	378	)	,
(	377	)	,
(	375	)	,
(	374	)	,
(	373	)	,
(	372	)	,
(	370	)	,
(	369	)	,
(	368	)	,
(	367	)	,
(	365	)	,
(	364	)	,
(	363	)	,
(	362	)	,
(	361	)	,
(	359	)	,
(	358	)	,
(	357	)	,
(	356	)	,
(	354	)	,
(	353	)	,
(	352	)	,
(	351	)	,
(	349	)	,
(	348	)	,
(	347	)	,
(	346	)	,
(	344	)	,
(	343	)	,
(	342	)	,
(	341	)	,
(	340	)	,
(	338	)	,
(	337	)	,
(	336	)	,
(	335	)	,
(	333	)	,
(	332	)	,
(	331	)	,
(	330	)	,
(	328	)	,
(	327	)	,
(	326	)	,
(	325	)	,
(	323	)	,
(	322	)	,
(	321	)	,
(	320	)	,
(	319	)	,
(	317	)	,
(	316	)	,
(	315	)	,
(	314	)	,
(	312	)	,
(	311	)	,
(	310	)	,
(	309	)	,
(	307	)	,
(	306	)	,
(	305	)	,
(	304	)	,
(	303	)	,
(	301	)	,
(	300	)	,
(	299	)	,
(	298	)	,
(	296	)	,
(	295	)	,
(	294	)	,
(	293	)	,
(	291	)	,
(	290	)	,
(	289	)	,
(	288	)	,
(	286	)	,
(	285	)	,
(	284	)	,
(	283	)	,
(	282	)	,
(	280	)	,
(	279	)	,
(	278	)	,
(	277	)	,
(	275	)	,
(	274	)	,
(	273	)	,
(	272	)	,
(	270	)	,
(	269	)	,
(	268	)	,
(	267	)	,
(	265	)	,
(	264	)	,
(	263	)	,
(	262	)	,
(	261	)	,
(	259	)	,
(	258	)	,
(	257	)	,
(	256	)	,
(	254	)	,
(	253	)	,
(	252	)	,
(	251	)	,
(	249	)	,
(	248	)	,
(	247	)	,
(	246	)	,
(	245	)	,
(	243	)	,
(	242	)	,
(	241	)	,
(	240	)	,
(	238	)	,
(	237	)	,
(	236	)	,
(	235	)	,
(	233	)	,
(	232	)	,
(	231	)	,
(	230	)	,
(	228	)	,
(	227	)	,
(	226	)	,
(	225	)	,
(	224	)	,
(	222	)	,
(	221	)	,
(	220	)	,
(	219	)	,
(	217	)	,
(	216	)	,
(	215	)	,
(	214	)	,
(	212	)	,
(	211	)	,
(	210	)	,
(	209	)	,
(	207	)	,
(	206	)	,
(	205	)	,
(	204	)	,
(	203	)	,
(	201	)	,
(	200	)	,
(	199	)	,
(	198	)	,
(	196	)	,
(	195	)	,
(	194	)	,
(	193	)	,
(	191	)	,
(	190	)	,
(	189	)	,
(	188	)	,
(	187	)	,
(	185	)	,
(	184	)	,
(	183	)	,
(	182	)	,
(	180	)	,
(	179	)	,
(	178	)	,
(	177	)	,
(	175	)	,
(	174	)	,
(	173	)	,
(	172	)	,
(	170	)	,
(	169	)	,
(	168	)	,
(	167	)	,
(	166	)	,
(	164	)	,
(	163	)	,
(	162	)	,
(	161	)	,
(	159	)	,
(	158	)	,
(	157	)	,
(	156	)	,
(	154	)	,
(	153	)	,
(	152	)	,
(	151	)	,
(	149	)	,
(	148	)	,
(	147	)	,
(	146	)	,
(	145	)	,
(	143	)	,
(	142	)	,
(	141	)	,
(	140	)	,
(	138	)	,
(	137	)	,
(	136	)	,
(	135	)	,
(	133	)	,
(	132	)	,
(	131	)	,
(	130	)	,
(	129	)	,
(	127	)	,
(	126	)	,
(	125	)	,
(	124	)	,
(	122	)	,
(	121	)	,
(	120	)	,
(	119	)	,
(	117	)	,
(	116	)	,
(	115	)	,
(	114	)	,
(	112	)	,
(	111	)	,
(	110	)	,
(	109	)	,
(	108	)	,
(	106	)	,
(	105	)	,
(	104	)	,
(	103	)	,
(	101	)	,
(	100	)	,
(	99	)	,
(	98	)	,
(	96	)	,
(	95	)	,
(	94	)	,
(	93	)	,
(	91	)	,
(	90	)	,
(	89	)	,
(	88	)	,
(	87	)	,
(	85	)	,
(	84	)	,
(	83	)	,
(	82	)	,
(	80	)	,
(	79	)	,
(	78	)	,
(	77	)	,
(	75	)	,
(	74	)	,
(	73	)	,
(	72	)	,
(	71	)	,
(	69	)	,
(	68	)	,
(	67	)	,
(	66	)	,
(	64	)	,
(	63	)	,
(	62	)	,
(	61	)	,
(	59	)	,
(	58	)	,
(	57	)	,
(	56	)	,
(	54	)	,
(	53	)	,
(	52	)	,
(	51	)	,
(	50	)	,
(	48	)	,
(	47	)	,
(	46	)	,
(	45	)	,
(	43	)	,
(	42	)	,
(	41	)	,
(	40	)	,
(	38	)	,
(	37	)	,
(	36	)	,
(	35	)	,
(	33	)	,
(	32	)	,
(	31	)	,
(	30	)	,
(	29	)	,
(	27	)	,
(	26	)	,
(	25	)	,
(	24	)	,
(	22	)	,
(	21	)	,
(	20	)	,
(	19	)	,
(	17	)	,
(	16	)	,
(	15	)	,
(	14	)	,
(	13	)	,
(	11	)	,
(	10	)	,
(	9	)	,
(	8	)	,
(	6	)	,
(	5	)	,
(	4	)	,
(	3	)	,
(	1	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)    -- array index 4095 (voltage = "111111111111" or 4095 mV), distance output 3787 (37.87 cm)

);


end package LUT_pkg;
