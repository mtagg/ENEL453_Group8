--file init for freeze entity