--test bench file init for freeze module