--only modifications to PWN_DAC were the enable functionality, reference the commented lines within the file for more info

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_PWM_DAC is
end entity;


--Apparently we dont need this for the demo